module delta_tb;

logic resetn = 1;
logic [2:0] delta = 0;
logic clk = 0;
logic [3:0] count;

initial begin
count = 0;
end

initial forever #10 clk = ~clk;

initial begin
delta = 3;
#240 delta = 2;
#200 delta = 7;
#900 delta = 0;
#2000 $stop;
end

initial begin
 #5 resetn = ~resetn;
 #5 resetn = ~resetn;
 #1760 resetn = ~resetn;
 #5 resetn = ~resetn;
end

initial forever #20 $strobe("counter value %d, delta value %d", count, delta);

delta uut_inst(.delta(delta), .count(count),.clk(clk), .resetn(resetn));

endmodule
